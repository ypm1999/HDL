`include "defines.v"

module IF (
	input wire 				clk,
	input wire 				rst,
	input wire 				rdy,

	input wire 				use_npc,
	input wire[31:0]		npc_addr,
	input wire[31:0]		ram_inst,
	input wire 				ram_inst_busy,
	input wire[4:0] 		stall,

	output reg[31:0] 		pc,
	output reg[31:0]		inst,
	output reg 				ram_inst_re,
	output reg[31:0]		ram_inst_addr,

	output reg 				stall_req
	);
	reg 		bj_stall, try_stall, rst_stall;

	always @ ( posedge clk ) begin
		if (rst == `RstEnable)begin
			pc <= -4;
			ram_inst_re <= `False_v;
			ram_inst_addr <= 32'hffffffff;
			try_stall <= `False_v;
			bj_stall <= `False_v;
		end
		else if(rdy == `True_v) begin
			if (stall[0] == `False_v) begin
				if (inst[6:4] == 3'b110 && !bj_stall)begin
					ram_inst_re <= `False_v;
					bj_stall <= `True_v;
				end
				else if (use_npc) begin
					pc <= npc_addr;
					ram_inst_re <= `True_v;
					ram_inst_addr <= npc_addr;
					try_stall <= ~try_stall;
					bj_stall <= `False_v;
				end
				else begin
					pc <= pc + 4;
					ram_inst_re <= `True_v;
					ram_inst_addr <= pc + 4;
					try_stall <= ~try_stall;
					bj_stall <= `False_v;
				end
			end
		end
	end

	always @ ( rst or ram_inst_busy ) begin
			if (rst) begin
				rst_stall <= `False_v;
				inst <= `ZeroWord;
			end
			else if(rdy == `True_v) begin
				if (ram_inst_re & !ram_inst_busy)begin
					rst_stall <= ~rst_stall;
					inst <= ram_inst;
				end
				else begin
					inst <= `ZeroWord;
				end
			end
		end

		always @ ( * ) begin
			if (rst)
				stall_req <= `False_v;
			else if (rdy) begin
				stall_req <= (try_stall ^ rst_stall);
			end
		end

endmodule // pc_reg
