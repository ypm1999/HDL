`include "defines.v"

module Ctrl (
	input wire 				clk,
	input wire 				rst,
	input wire 				rdy,

	input wire 				if_stall,
	input wire 				ex_stall,
	input wire 				if_stall,
	input wire 				if_stall,
	);

endmodule // Ctrl
