`include "defines.v"

module MemoryCtrl (

	);

endmodule // MemoryCtrl
